magic
tech scmos
timestamp 1732295240
<< nwell >>
rect -45 -6 1913 14
<< ntransistor >>
rect -29 -64 -27 -60
rect 7 -64 9 -60
rect 49 -64 51 -60
rect 67 -64 69 -60
rect 97 -64 99 -60
rect 132 -64 134 -60
rect 150 -64 152 -60
rect 180 -64 182 -60
rect 215 -64 217 -60
rect 233 -64 235 -60
rect 263 -64 265 -60
rect 298 -64 300 -60
rect 316 -64 318 -60
rect 346 -64 348 -60
rect 399 -64 401 -60
rect 417 -64 419 -60
rect 447 -64 449 -60
rect 496 -64 498 -60
rect 514 -64 516 -60
rect 562 -64 564 -60
rect 619 -64 621 -60
rect 655 -64 657 -60
rect 697 -64 699 -60
rect 715 -64 717 -60
rect 745 -64 747 -60
rect 780 -64 782 -60
rect 798 -64 800 -60
rect 828 -64 830 -60
rect 863 -64 865 -60
rect 881 -64 883 -60
rect 911 -64 913 -60
rect 954 -64 956 -60
rect 990 -64 992 -60
rect 1032 -64 1034 -60
rect 1050 -64 1052 -60
rect 1080 -64 1082 -60
rect 1115 -64 1117 -60
rect 1133 -64 1135 -60
rect 1163 -64 1165 -60
rect 1198 -64 1200 -60
rect 1216 -64 1218 -60
rect 1246 -64 1248 -60
rect 1281 -64 1283 -60
rect 1299 -64 1301 -60
rect 1329 -64 1331 -60
rect 1382 -64 1384 -60
rect 1400 -64 1402 -60
rect 1430 -64 1432 -60
rect 1479 -64 1481 -60
rect 1497 -64 1499 -60
rect 1545 -64 1547 -60
rect 1602 -64 1604 -60
rect 1638 -64 1640 -60
rect 1680 -64 1682 -60
rect 1698 -64 1700 -60
rect 1728 -64 1730 -60
rect 1763 -64 1765 -60
rect 1781 -64 1783 -60
rect 1811 -64 1813 -60
rect 1846 -64 1848 -60
rect 1864 -64 1866 -60
rect 1894 -64 1896 -60
<< ptransistor >>
rect -29 0 -27 8
rect 7 0 9 8
rect 49 0 51 8
rect 67 0 69 8
rect 97 0 99 8
rect 132 0 134 8
rect 150 0 152 8
rect 180 0 182 8
rect 215 0 217 8
rect 233 0 235 8
rect 263 0 265 8
rect 298 0 300 8
rect 316 0 318 8
rect 346 0 348 8
rect 399 0 401 8
rect 417 0 419 8
rect 447 0 449 8
rect 496 0 498 8
rect 514 0 516 8
rect 562 0 564 8
rect 619 0 621 8
rect 655 0 657 8
rect 697 0 699 8
rect 715 0 717 8
rect 745 0 747 8
rect 780 0 782 8
rect 798 0 800 8
rect 828 0 830 8
rect 863 0 865 8
rect 881 0 883 8
rect 911 0 913 8
rect 954 0 956 8
rect 990 0 992 8
rect 1032 0 1034 8
rect 1050 0 1052 8
rect 1080 0 1082 8
rect 1115 0 1117 8
rect 1133 0 1135 8
rect 1163 0 1165 8
rect 1198 0 1200 8
rect 1216 0 1218 8
rect 1246 0 1248 8
rect 1281 0 1283 8
rect 1299 0 1301 8
rect 1329 0 1331 8
rect 1382 0 1384 8
rect 1400 0 1402 8
rect 1430 0 1432 8
rect 1479 0 1481 8
rect 1497 0 1499 8
rect 1545 0 1547 8
rect 1602 0 1604 8
rect 1638 0 1640 8
rect 1680 0 1682 8
rect 1698 0 1700 8
rect 1728 0 1730 8
rect 1763 0 1765 8
rect 1781 0 1783 8
rect 1811 0 1813 8
rect 1846 0 1848 8
rect 1864 0 1866 8
rect 1894 0 1896 8
<< ndiffusion >>
rect -35 -64 -29 -60
rect -27 -64 -21 -60
rect 1 -64 7 -60
rect 9 -64 15 -60
rect 43 -64 49 -60
rect 51 -64 67 -60
rect 69 -64 71 -60
rect 91 -64 97 -60
rect 99 -64 105 -60
rect 126 -64 132 -60
rect 134 -64 150 -60
rect 152 -64 154 -60
rect 174 -64 180 -60
rect 182 -64 188 -60
rect 209 -64 215 -60
rect 217 -64 219 -60
rect 223 -64 233 -60
rect 235 -64 237 -60
rect 257 -64 263 -60
rect 265 -64 271 -60
rect 292 -64 298 -60
rect 300 -64 316 -60
rect 318 -64 320 -60
rect 340 -64 346 -60
rect 348 -64 354 -60
rect 393 -64 399 -60
rect 401 -64 417 -60
rect 419 -64 421 -60
rect 441 -64 447 -60
rect 449 -64 455 -60
rect 490 -64 496 -60
rect 498 -64 500 -60
rect 504 -64 514 -60
rect 516 -64 518 -60
rect 556 -64 562 -60
rect 564 -64 570 -60
rect 613 -64 619 -60
rect 621 -64 627 -60
rect 649 -64 655 -60
rect 657 -64 663 -60
rect 691 -64 697 -60
rect 699 -64 715 -60
rect 717 -64 719 -60
rect 739 -64 745 -60
rect 747 -64 753 -60
rect 774 -64 780 -60
rect 782 -64 798 -60
rect 800 -64 802 -60
rect 822 -64 828 -60
rect 830 -64 836 -60
rect 857 -64 863 -60
rect 865 -64 867 -60
rect 871 -64 881 -60
rect 883 -64 885 -60
rect 905 -64 911 -60
rect 913 -64 919 -60
rect 948 -64 954 -60
rect 956 -64 962 -60
rect 984 -64 990 -60
rect 992 -64 998 -60
rect 1026 -64 1032 -60
rect 1034 -64 1050 -60
rect 1052 -64 1054 -60
rect 1074 -64 1080 -60
rect 1082 -64 1088 -60
rect 1109 -64 1115 -60
rect 1117 -64 1133 -60
rect 1135 -64 1137 -60
rect 1157 -64 1163 -60
rect 1165 -64 1171 -60
rect 1192 -64 1198 -60
rect 1200 -64 1202 -60
rect 1206 -64 1216 -60
rect 1218 -64 1220 -60
rect 1240 -64 1246 -60
rect 1248 -64 1254 -60
rect 1275 -64 1281 -60
rect 1283 -64 1299 -60
rect 1301 -64 1303 -60
rect 1323 -64 1329 -60
rect 1331 -64 1337 -60
rect 1376 -64 1382 -60
rect 1384 -64 1400 -60
rect 1402 -64 1404 -60
rect 1424 -64 1430 -60
rect 1432 -64 1438 -60
rect 1473 -64 1479 -60
rect 1481 -64 1483 -60
rect 1487 -64 1497 -60
rect 1499 -64 1501 -60
rect 1539 -64 1545 -60
rect 1547 -64 1553 -60
rect 1596 -64 1602 -60
rect 1604 -64 1610 -60
rect 1632 -64 1638 -60
rect 1640 -64 1646 -60
rect 1674 -64 1680 -60
rect 1682 -64 1698 -60
rect 1700 -64 1702 -60
rect 1722 -64 1728 -60
rect 1730 -64 1736 -60
rect 1757 -64 1763 -60
rect 1765 -64 1781 -60
rect 1783 -64 1785 -60
rect 1805 -64 1811 -60
rect 1813 -64 1819 -60
rect 1840 -64 1846 -60
rect 1848 -64 1850 -60
rect 1854 -64 1864 -60
rect 1866 -64 1868 -60
rect 1888 -64 1894 -60
rect 1896 -64 1902 -60
<< pdiffusion >>
rect -35 0 -29 8
rect -27 0 -21 8
rect 1 0 7 8
rect 9 0 15 8
rect 43 0 49 8
rect 51 0 53 8
rect 57 0 67 8
rect 69 0 71 8
rect 91 0 97 8
rect 99 0 105 8
rect 126 0 132 8
rect 134 0 136 8
rect 140 0 150 8
rect 152 0 154 8
rect 174 0 180 8
rect 182 0 188 8
rect 209 0 215 8
rect 217 0 233 8
rect 235 0 237 8
rect 257 0 263 8
rect 265 0 271 8
rect 292 0 298 8
rect 300 0 302 8
rect 306 0 316 8
rect 318 0 320 8
rect 340 0 346 8
rect 348 0 354 8
rect 393 0 399 8
rect 401 0 403 8
rect 407 0 417 8
rect 419 0 421 8
rect 441 0 447 8
rect 449 0 455 8
rect 490 0 496 8
rect 498 0 514 8
rect 516 0 518 8
rect 556 0 562 8
rect 564 0 570 8
rect 613 0 619 8
rect 621 0 627 8
rect 649 0 655 8
rect 657 0 663 8
rect 691 0 697 8
rect 699 0 701 8
rect 705 0 715 8
rect 717 0 719 8
rect 739 0 745 8
rect 747 0 753 8
rect 774 0 780 8
rect 782 0 784 8
rect 788 0 798 8
rect 800 0 802 8
rect 822 0 828 8
rect 830 0 836 8
rect 857 0 863 8
rect 865 0 881 8
rect 883 0 885 8
rect 905 0 911 8
rect 913 0 919 8
rect 948 0 954 8
rect 956 0 962 8
rect 984 0 990 8
rect 992 0 998 8
rect 1026 0 1032 8
rect 1034 0 1036 8
rect 1040 0 1050 8
rect 1052 0 1054 8
rect 1074 0 1080 8
rect 1082 0 1088 8
rect 1109 0 1115 8
rect 1117 0 1119 8
rect 1123 0 1133 8
rect 1135 0 1137 8
rect 1157 0 1163 8
rect 1165 0 1171 8
rect 1192 0 1198 8
rect 1200 0 1216 8
rect 1218 0 1220 8
rect 1240 0 1246 8
rect 1248 0 1254 8
rect 1275 0 1281 8
rect 1283 0 1285 8
rect 1289 0 1299 8
rect 1301 0 1303 8
rect 1323 0 1329 8
rect 1331 0 1337 8
rect 1376 0 1382 8
rect 1384 0 1386 8
rect 1390 0 1400 8
rect 1402 0 1404 8
rect 1424 0 1430 8
rect 1432 0 1438 8
rect 1473 0 1479 8
rect 1481 0 1497 8
rect 1499 0 1501 8
rect 1539 0 1545 8
rect 1547 0 1553 8
rect 1596 0 1602 8
rect 1604 0 1610 8
rect 1632 0 1638 8
rect 1640 0 1646 8
rect 1674 0 1680 8
rect 1682 0 1684 8
rect 1688 0 1698 8
rect 1700 0 1702 8
rect 1722 0 1728 8
rect 1730 0 1736 8
rect 1757 0 1763 8
rect 1765 0 1767 8
rect 1771 0 1781 8
rect 1783 0 1785 8
rect 1805 0 1811 8
rect 1813 0 1819 8
rect 1840 0 1846 8
rect 1848 0 1864 8
rect 1866 0 1868 8
rect 1888 0 1894 8
rect 1896 0 1902 8
<< ndcontact >>
rect -39 -64 -35 -60
rect -21 -64 -17 -60
rect -3 -64 1 -60
rect 15 -64 19 -60
rect 39 -64 43 -60
rect 71 -64 75 -60
rect 87 -64 91 -60
rect 105 -64 109 -60
rect 122 -64 126 -60
rect 154 -64 158 -60
rect 170 -64 174 -60
rect 188 -64 192 -60
rect 205 -64 209 -60
rect 219 -64 223 -60
rect 237 -64 241 -60
rect 253 -64 257 -60
rect 271 -64 275 -60
rect 288 -64 292 -60
rect 320 -64 324 -60
rect 336 -64 340 -60
rect 354 -64 358 -60
rect 389 -64 393 -60
rect 421 -64 425 -60
rect 437 -64 441 -60
rect 455 -64 459 -60
rect 486 -64 490 -60
rect 500 -64 504 -60
rect 518 -64 522 -60
rect 552 -64 556 -60
rect 570 -64 574 -60
rect 609 -64 613 -60
rect 627 -64 631 -60
rect 645 -64 649 -60
rect 663 -64 667 -60
rect 687 -64 691 -60
rect 719 -64 723 -60
rect 735 -64 739 -60
rect 753 -64 757 -60
rect 770 -64 774 -60
rect 802 -64 806 -60
rect 818 -64 822 -60
rect 836 -64 840 -60
rect 853 -64 857 -60
rect 867 -64 871 -60
rect 885 -64 889 -60
rect 901 -64 905 -60
rect 919 -64 923 -60
rect 944 -64 948 -60
rect 962 -64 966 -60
rect 980 -64 984 -60
rect 998 -64 1002 -60
rect 1022 -64 1026 -60
rect 1054 -64 1058 -60
rect 1070 -64 1074 -60
rect 1088 -64 1092 -60
rect 1105 -64 1109 -60
rect 1137 -64 1141 -60
rect 1153 -64 1157 -60
rect 1171 -64 1175 -60
rect 1188 -64 1192 -60
rect 1202 -64 1206 -60
rect 1220 -64 1224 -60
rect 1236 -64 1240 -60
rect 1254 -64 1258 -60
rect 1271 -64 1275 -60
rect 1303 -64 1307 -60
rect 1319 -64 1323 -60
rect 1337 -64 1341 -60
rect 1372 -64 1376 -60
rect 1404 -64 1408 -60
rect 1420 -64 1424 -60
rect 1438 -64 1442 -60
rect 1469 -64 1473 -60
rect 1483 -64 1487 -60
rect 1501 -64 1505 -60
rect 1535 -64 1539 -60
rect 1553 -64 1557 -60
rect 1592 -64 1596 -60
rect 1610 -64 1614 -60
rect 1628 -64 1632 -60
rect 1646 -64 1650 -60
rect 1670 -64 1674 -60
rect 1702 -64 1706 -60
rect 1718 -64 1722 -60
rect 1736 -64 1740 -60
rect 1753 -64 1757 -60
rect 1785 -64 1789 -60
rect 1801 -64 1805 -60
rect 1819 -64 1823 -60
rect 1836 -64 1840 -60
rect 1850 -64 1854 -60
rect 1868 -64 1872 -60
rect 1884 -64 1888 -60
rect 1902 -64 1906 -60
<< pdcontact >>
rect -39 0 -35 8
rect -21 0 -17 8
rect -3 0 1 8
rect 15 0 19 8
rect 39 0 43 8
rect 53 0 57 8
rect 71 0 75 8
rect 87 0 91 8
rect 105 0 109 8
rect 122 0 126 8
rect 136 0 140 8
rect 154 0 158 8
rect 170 0 174 8
rect 188 0 192 8
rect 205 0 209 8
rect 237 0 241 8
rect 253 0 257 8
rect 271 0 275 8
rect 288 0 292 8
rect 302 0 306 8
rect 320 0 324 8
rect 336 0 340 8
rect 354 0 358 8
rect 389 0 393 8
rect 403 0 407 8
rect 421 0 425 8
rect 437 0 441 8
rect 455 0 459 8
rect 486 0 490 8
rect 518 0 522 8
rect 552 0 556 8
rect 570 0 574 8
rect 609 0 613 8
rect 627 0 631 8
rect 645 0 649 8
rect 663 0 667 8
rect 687 0 691 8
rect 701 0 705 8
rect 719 0 723 8
rect 735 0 739 8
rect 753 0 757 8
rect 770 0 774 8
rect 784 0 788 8
rect 802 0 806 8
rect 818 0 822 8
rect 836 0 840 8
rect 853 0 857 8
rect 885 0 889 8
rect 901 0 905 8
rect 919 0 923 8
rect 944 0 948 8
rect 962 0 966 8
rect 980 0 984 8
rect 998 0 1002 8
rect 1022 0 1026 8
rect 1036 0 1040 8
rect 1054 0 1058 8
rect 1070 0 1074 8
rect 1088 0 1092 8
rect 1105 0 1109 8
rect 1119 0 1123 8
rect 1137 0 1141 8
rect 1153 0 1157 8
rect 1171 0 1175 8
rect 1188 0 1192 8
rect 1220 0 1224 8
rect 1236 0 1240 8
rect 1254 0 1258 8
rect 1271 0 1275 8
rect 1285 0 1289 8
rect 1303 0 1307 8
rect 1319 0 1323 8
rect 1337 0 1341 8
rect 1372 0 1376 8
rect 1386 0 1390 8
rect 1404 0 1408 8
rect 1420 0 1424 8
rect 1438 0 1442 8
rect 1469 0 1473 8
rect 1501 0 1505 8
rect 1535 0 1539 8
rect 1553 0 1557 8
rect 1592 0 1596 8
rect 1610 0 1614 8
rect 1628 0 1632 8
rect 1646 0 1650 8
rect 1670 0 1674 8
rect 1684 0 1688 8
rect 1702 0 1706 8
rect 1718 0 1722 8
rect 1736 0 1740 8
rect 1753 0 1757 8
rect 1767 0 1771 8
rect 1785 0 1789 8
rect 1801 0 1805 8
rect 1819 0 1823 8
rect 1836 0 1840 8
rect 1868 0 1872 8
rect 1884 0 1888 8
rect 1902 0 1906 8
<< psubstratepcontact >>
rect -39 -76 -35 -72
rect -25 -76 -21 -72
rect -14 -76 -10 -72
rect -3 -76 1 -72
rect 11 -76 15 -72
rect 22 -76 26 -72
rect 39 -76 43 -72
rect 53 -76 57 -72
rect 67 -76 71 -72
rect 87 -76 91 -72
rect 101 -76 105 -72
rect 112 -76 116 -72
rect 122 -76 126 -72
rect 136 -76 140 -72
rect 150 -76 154 -72
rect 170 -76 174 -72
rect 184 -76 188 -72
rect 195 -76 199 -72
rect 205 -76 209 -72
rect 219 -76 223 -72
rect 237 -76 241 -72
rect 253 -76 257 -72
rect 267 -76 271 -72
rect 278 -76 282 -72
rect 288 -76 292 -72
rect 302 -76 306 -72
rect 316 -76 320 -72
rect 336 -76 340 -72
rect 350 -76 354 -72
rect 361 -76 365 -72
rect 389 -76 393 -72
rect 403 -76 407 -72
rect 417 -76 421 -72
rect 437 -76 441 -72
rect 451 -76 455 -72
rect 462 -76 466 -72
rect 486 -76 490 -72
rect 500 -76 504 -72
rect 518 -76 522 -72
rect 552 -76 556 -72
rect 566 -76 570 -72
rect 577 -76 581 -72
rect 609 -76 613 -72
rect 623 -76 627 -72
rect 634 -76 638 -72
rect 645 -76 649 -72
rect 659 -76 663 -72
rect 670 -76 674 -72
rect 687 -76 691 -72
rect 701 -76 705 -72
rect 715 -76 719 -72
rect 735 -76 739 -72
rect 749 -76 753 -72
rect 760 -76 764 -72
rect 770 -76 774 -72
rect 784 -76 788 -72
rect 798 -76 802 -72
rect 818 -76 822 -72
rect 832 -76 836 -72
rect 843 -76 847 -72
rect 853 -76 857 -72
rect 867 -76 871 -72
rect 885 -76 889 -72
rect 901 -76 905 -72
rect 915 -76 919 -72
rect 926 -76 930 -72
rect 944 -76 948 -72
rect 958 -76 962 -72
rect 969 -76 973 -72
rect 980 -76 984 -72
rect 994 -76 998 -72
rect 1005 -76 1009 -72
rect 1022 -76 1026 -72
rect 1036 -76 1040 -72
rect 1050 -76 1054 -72
rect 1070 -76 1074 -72
rect 1084 -76 1088 -72
rect 1095 -76 1099 -72
rect 1105 -76 1109 -72
rect 1119 -76 1123 -72
rect 1133 -76 1137 -72
rect 1153 -76 1157 -72
rect 1167 -76 1171 -72
rect 1178 -76 1182 -72
rect 1188 -76 1192 -72
rect 1202 -76 1206 -72
rect 1220 -76 1224 -72
rect 1236 -76 1240 -72
rect 1250 -76 1254 -72
rect 1261 -76 1265 -72
rect 1271 -76 1275 -72
rect 1285 -76 1289 -72
rect 1299 -76 1303 -72
rect 1319 -76 1323 -72
rect 1333 -76 1337 -72
rect 1344 -76 1348 -72
rect 1372 -76 1376 -72
rect 1386 -76 1390 -72
rect 1400 -76 1404 -72
rect 1420 -76 1424 -72
rect 1434 -76 1438 -72
rect 1445 -76 1449 -72
rect 1469 -76 1473 -72
rect 1483 -76 1487 -72
rect 1501 -76 1505 -72
rect 1535 -76 1539 -72
rect 1549 -76 1553 -72
rect 1560 -76 1564 -72
rect 1592 -76 1596 -72
rect 1606 -76 1610 -72
rect 1617 -76 1621 -72
rect 1628 -76 1632 -72
rect 1642 -76 1646 -72
rect 1653 -76 1657 -72
rect 1670 -76 1674 -72
rect 1684 -76 1688 -72
rect 1698 -76 1702 -72
rect 1718 -76 1722 -72
rect 1732 -76 1736 -72
rect 1743 -76 1747 -72
rect 1753 -76 1757 -72
rect 1767 -76 1771 -72
rect 1781 -76 1785 -72
rect 1801 -76 1805 -72
rect 1815 -76 1819 -72
rect 1826 -76 1830 -72
rect 1836 -76 1840 -72
rect 1850 -76 1854 -72
rect 1868 -76 1872 -72
rect 1884 -76 1888 -72
rect 1898 -76 1902 -72
rect 1909 -76 1913 -72
<< nsubstratencontact >>
rect -39 20 -35 24
rect -28 20 -24 24
rect -17 20 -13 24
rect -3 20 1 24
rect 8 20 12 24
rect 19 20 23 24
rect 39 20 43 24
rect 53 20 57 24
rect 71 20 75 24
rect 87 20 91 24
rect 98 20 102 24
rect 109 20 113 24
rect 122 20 126 24
rect 136 20 140 24
rect 154 20 158 24
rect 170 20 174 24
rect 181 20 185 24
rect 192 20 196 24
rect 205 20 209 24
rect 219 20 223 24
rect 237 20 241 24
rect 253 20 257 24
rect 264 20 268 24
rect 275 20 279 24
rect 288 20 292 24
rect 302 20 306 24
rect 320 20 324 24
rect 336 20 340 24
rect 347 20 351 24
rect 358 20 362 24
rect 389 20 393 24
rect 403 20 407 24
rect 421 20 425 24
rect 437 20 441 24
rect 448 20 452 24
rect 459 20 463 24
rect 486 20 490 24
rect 500 20 504 24
rect 518 20 522 24
rect 552 20 556 24
rect 563 20 567 24
rect 574 20 578 24
rect 609 20 613 24
rect 620 20 624 24
rect 631 20 635 24
rect 645 20 649 24
rect 656 20 660 24
rect 667 20 671 24
rect 687 20 691 24
rect 701 20 705 24
rect 719 20 723 24
rect 735 20 739 24
rect 746 20 750 24
rect 757 20 761 24
rect 770 20 774 24
rect 784 20 788 24
rect 802 20 806 24
rect 818 20 822 24
rect 829 20 833 24
rect 840 20 844 24
rect 853 20 857 24
rect 867 20 871 24
rect 885 20 889 24
rect 901 20 905 24
rect 912 20 916 24
rect 923 20 927 24
rect 944 20 948 24
rect 955 20 959 24
rect 966 20 970 24
rect 980 20 984 24
rect 991 20 995 24
rect 1002 20 1006 24
rect 1022 20 1026 24
rect 1036 20 1040 24
rect 1054 20 1058 24
rect 1070 20 1074 24
rect 1081 20 1085 24
rect 1092 20 1096 24
rect 1105 20 1109 24
rect 1119 20 1123 24
rect 1137 20 1141 24
rect 1153 20 1157 24
rect 1164 20 1168 24
rect 1175 20 1179 24
rect 1188 20 1192 24
rect 1202 20 1206 24
rect 1220 20 1224 24
rect 1236 20 1240 24
rect 1247 20 1251 24
rect 1258 20 1262 24
rect 1271 20 1275 24
rect 1285 20 1289 24
rect 1303 20 1307 24
rect 1319 20 1323 24
rect 1330 20 1334 24
rect 1341 20 1345 24
rect 1372 20 1376 24
rect 1386 20 1390 24
rect 1404 20 1408 24
rect 1420 20 1424 24
rect 1431 20 1435 24
rect 1442 20 1446 24
rect 1469 20 1473 24
rect 1483 20 1487 24
rect 1501 20 1505 24
rect 1535 20 1539 24
rect 1546 20 1550 24
rect 1557 20 1561 24
rect 1592 20 1596 24
rect 1603 20 1607 24
rect 1614 20 1618 24
rect 1628 20 1632 24
rect 1639 20 1643 24
rect 1650 20 1654 24
rect 1670 20 1674 24
rect 1684 20 1688 24
rect 1702 20 1706 24
rect 1718 20 1722 24
rect 1729 20 1733 24
rect 1740 20 1744 24
rect 1753 20 1757 24
rect 1767 20 1771 24
rect 1785 20 1789 24
rect 1801 20 1805 24
rect 1812 20 1816 24
rect 1823 20 1827 24
rect 1836 20 1840 24
rect 1850 20 1854 24
rect 1868 20 1872 24
rect 1884 20 1888 24
rect 1895 20 1899 24
rect 1906 20 1910 24
<< polysilicon >>
rect -29 8 -27 12
rect 7 8 9 12
rect 49 8 51 12
rect 67 8 69 12
rect 97 8 99 12
rect 132 8 134 12
rect 150 8 152 12
rect 180 8 182 12
rect 215 8 217 12
rect 233 8 235 12
rect 263 8 265 12
rect 298 8 300 12
rect 316 8 318 12
rect 346 8 348 12
rect 399 8 401 12
rect 417 8 419 12
rect 447 8 449 12
rect 496 8 498 12
rect 514 8 516 12
rect 562 8 564 12
rect 619 8 621 12
rect 655 8 657 12
rect 697 8 699 12
rect 715 8 717 12
rect 745 8 747 12
rect 780 8 782 12
rect 798 8 800 12
rect 828 8 830 12
rect 863 8 865 12
rect 881 8 883 12
rect 911 8 913 12
rect 954 8 956 12
rect 990 8 992 12
rect 1032 8 1034 12
rect 1050 8 1052 12
rect 1080 8 1082 12
rect 1115 8 1117 12
rect 1133 8 1135 12
rect 1163 8 1165 12
rect 1198 8 1200 12
rect 1216 8 1218 12
rect 1246 8 1248 12
rect 1281 8 1283 12
rect 1299 8 1301 12
rect 1329 8 1331 12
rect 1382 8 1384 12
rect 1400 8 1402 12
rect 1430 8 1432 12
rect 1479 8 1481 12
rect 1497 8 1499 12
rect 1545 8 1547 12
rect 1602 8 1604 12
rect 1638 8 1640 12
rect 1680 8 1682 12
rect 1698 8 1700 12
rect 1728 8 1730 12
rect 1763 8 1765 12
rect 1781 8 1783 12
rect 1811 8 1813 12
rect 1846 8 1848 12
rect 1864 8 1866 12
rect 1894 8 1896 12
rect -29 -31 -27 0
rect 7 -31 9 0
rect 49 -15 51 0
rect 50 -19 51 -15
rect -28 -35 -27 -31
rect 8 -35 9 -31
rect -29 -60 -27 -35
rect 7 -60 9 -35
rect 49 -60 51 -19
rect 67 -43 69 0
rect 97 -32 99 0
rect 132 -14 134 0
rect 133 -18 134 -14
rect 98 -36 99 -32
rect 68 -47 69 -43
rect 67 -60 69 -47
rect 97 -60 99 -36
rect 132 -60 134 -18
rect 150 -43 152 0
rect 180 -32 182 0
rect 215 -32 217 0
rect 233 -15 235 0
rect 234 -19 235 -15
rect 181 -36 182 -32
rect 216 -36 217 -32
rect 151 -47 152 -43
rect 150 -60 152 -47
rect 180 -60 182 -36
rect 215 -60 217 -36
rect 233 -60 235 -19
rect 263 -32 265 0
rect 298 -7 300 0
rect 299 -11 300 -7
rect 264 -36 265 -32
rect 263 -60 265 -36
rect 298 -60 300 -11
rect 316 -43 318 0
rect 346 -32 348 0
rect 399 -11 401 0
rect 400 -15 401 -11
rect 347 -36 348 -32
rect 317 -47 318 -43
rect 316 -60 318 -47
rect 346 -60 348 -36
rect 399 -60 401 -15
rect 417 -33 419 0
rect 447 -26 449 0
rect 448 -30 449 -26
rect 418 -37 419 -33
rect 417 -60 419 -37
rect 447 -60 449 -30
rect 496 -34 498 0
rect 514 -11 516 0
rect 515 -15 516 -11
rect 497 -38 498 -34
rect 496 -60 498 -38
rect 514 -60 516 -15
rect 562 -32 564 0
rect 619 -31 621 0
rect 655 -31 657 0
rect 697 -15 699 0
rect 698 -19 699 -15
rect 563 -36 564 -32
rect 620 -35 621 -31
rect 656 -35 657 -31
rect 562 -60 564 -36
rect 619 -60 621 -35
rect 655 -60 657 -35
rect 697 -60 699 -19
rect 715 -43 717 0
rect 745 -32 747 0
rect 780 -14 782 0
rect 781 -18 782 -14
rect 746 -36 747 -32
rect 716 -47 717 -43
rect 715 -60 717 -47
rect 745 -60 747 -36
rect 780 -60 782 -18
rect 798 -43 800 0
rect 828 -32 830 0
rect 863 -32 865 0
rect 881 -15 883 0
rect 882 -19 883 -15
rect 829 -36 830 -32
rect 864 -36 865 -32
rect 799 -47 800 -43
rect 798 -60 800 -47
rect 828 -60 830 -36
rect 863 -60 865 -36
rect 881 -60 883 -19
rect 911 -32 913 0
rect 954 -31 956 0
rect 990 -31 992 0
rect 1032 -15 1034 0
rect 1033 -19 1034 -15
rect 912 -36 913 -32
rect 955 -35 956 -31
rect 991 -35 992 -31
rect 911 -60 913 -36
rect 954 -60 956 -35
rect 990 -60 992 -35
rect 1032 -60 1034 -19
rect 1050 -43 1052 0
rect 1080 -32 1082 0
rect 1115 -14 1117 0
rect 1116 -18 1117 -14
rect 1081 -36 1082 -32
rect 1051 -47 1052 -43
rect 1050 -60 1052 -47
rect 1080 -60 1082 -36
rect 1115 -60 1117 -18
rect 1133 -43 1135 0
rect 1163 -32 1165 0
rect 1198 -32 1200 0
rect 1216 -15 1218 0
rect 1217 -19 1218 -15
rect 1164 -36 1165 -32
rect 1199 -36 1200 -32
rect 1134 -47 1135 -43
rect 1133 -60 1135 -47
rect 1163 -60 1165 -36
rect 1198 -60 1200 -36
rect 1216 -60 1218 -19
rect 1246 -32 1248 0
rect 1281 -7 1283 0
rect 1282 -11 1283 -7
rect 1247 -36 1248 -32
rect 1246 -60 1248 -36
rect 1281 -60 1283 -11
rect 1299 -43 1301 0
rect 1329 -32 1331 0
rect 1382 -11 1384 0
rect 1383 -15 1384 -11
rect 1330 -36 1331 -32
rect 1300 -47 1301 -43
rect 1299 -60 1301 -47
rect 1329 -60 1331 -36
rect 1382 -60 1384 -15
rect 1400 -33 1402 0
rect 1430 -26 1432 0
rect 1431 -30 1432 -26
rect 1401 -37 1402 -33
rect 1400 -60 1402 -37
rect 1430 -60 1432 -30
rect 1479 -34 1481 0
rect 1497 -11 1499 0
rect 1498 -15 1499 -11
rect 1480 -38 1481 -34
rect 1479 -60 1481 -38
rect 1497 -60 1499 -15
rect 1545 -32 1547 0
rect 1602 -31 1604 0
rect 1638 -31 1640 0
rect 1680 -15 1682 0
rect 1681 -19 1682 -15
rect 1546 -36 1547 -32
rect 1603 -35 1604 -31
rect 1639 -35 1640 -31
rect 1545 -60 1547 -36
rect 1602 -60 1604 -35
rect 1638 -60 1640 -35
rect 1680 -60 1682 -19
rect 1698 -43 1700 0
rect 1728 -32 1730 0
rect 1763 -14 1765 0
rect 1764 -18 1765 -14
rect 1729 -36 1730 -32
rect 1699 -47 1700 -43
rect 1698 -60 1700 -47
rect 1728 -60 1730 -36
rect 1763 -60 1765 -18
rect 1781 -43 1783 0
rect 1811 -32 1813 0
rect 1846 -32 1848 0
rect 1864 -15 1866 0
rect 1865 -19 1866 -15
rect 1812 -36 1813 -32
rect 1847 -36 1848 -32
rect 1782 -47 1783 -43
rect 1781 -60 1783 -47
rect 1811 -60 1813 -36
rect 1846 -60 1848 -36
rect 1864 -60 1866 -19
rect 1894 -32 1896 0
rect 1895 -36 1896 -32
rect 1894 -60 1896 -36
rect -29 -67 -27 -64
rect 7 -67 9 -64
rect 49 -67 51 -64
rect 67 -68 69 -64
rect 97 -67 99 -64
rect 132 -67 134 -64
rect 150 -68 152 -64
rect 180 -67 182 -64
rect 215 -67 217 -64
rect 233 -68 235 -64
rect 263 -67 265 -64
rect 298 -67 300 -64
rect 316 -68 318 -64
rect 346 -67 348 -64
rect 399 -67 401 -64
rect 417 -68 419 -64
rect 447 -67 449 -64
rect 496 -67 498 -64
rect 514 -68 516 -64
rect 562 -67 564 -64
rect 619 -67 621 -64
rect 655 -67 657 -64
rect 697 -67 699 -64
rect 715 -68 717 -64
rect 745 -67 747 -64
rect 780 -67 782 -64
rect 798 -68 800 -64
rect 828 -67 830 -64
rect 863 -67 865 -64
rect 881 -68 883 -64
rect 911 -67 913 -64
rect 954 -67 956 -64
rect 990 -67 992 -64
rect 1032 -67 1034 -64
rect 1050 -68 1052 -64
rect 1080 -67 1082 -64
rect 1115 -67 1117 -64
rect 1133 -68 1135 -64
rect 1163 -67 1165 -64
rect 1198 -67 1200 -64
rect 1216 -68 1218 -64
rect 1246 -67 1248 -64
rect 1281 -67 1283 -64
rect 1299 -68 1301 -64
rect 1329 -67 1331 -64
rect 1382 -67 1384 -64
rect 1400 -68 1402 -64
rect 1430 -67 1432 -64
rect 1479 -67 1481 -64
rect 1497 -68 1499 -64
rect 1545 -67 1547 -64
rect 1602 -67 1604 -64
rect 1638 -67 1640 -64
rect 1680 -67 1682 -64
rect 1698 -68 1700 -64
rect 1728 -67 1730 -64
rect 1763 -67 1765 -64
rect 1781 -68 1783 -64
rect 1811 -67 1813 -64
rect 1846 -67 1848 -64
rect 1864 -68 1866 -64
rect 1894 -67 1896 -64
<< polycontact >>
rect 46 -19 50 -15
rect -32 -35 -28 -31
rect 4 -35 8 -31
rect 129 -18 133 -14
rect 94 -36 98 -32
rect 64 -47 68 -43
rect 230 -19 234 -15
rect 177 -36 181 -32
rect 212 -36 216 -32
rect 147 -47 151 -43
rect 295 -11 299 -7
rect 260 -36 264 -32
rect 396 -15 400 -11
rect 343 -36 347 -32
rect 313 -47 317 -43
rect 444 -30 448 -26
rect 414 -37 418 -33
rect 511 -15 515 -11
rect 493 -38 497 -34
rect 694 -19 698 -15
rect 559 -36 563 -32
rect 616 -35 620 -31
rect 652 -35 656 -31
rect 777 -18 781 -14
rect 742 -36 746 -32
rect 712 -47 716 -43
rect 878 -19 882 -15
rect 825 -36 829 -32
rect 860 -36 864 -32
rect 795 -47 799 -43
rect 1029 -19 1033 -15
rect 908 -36 912 -32
rect 951 -35 955 -31
rect 987 -35 991 -31
rect 1112 -18 1116 -14
rect 1077 -36 1081 -32
rect 1047 -47 1051 -43
rect 1213 -19 1217 -15
rect 1160 -36 1164 -32
rect 1195 -36 1199 -32
rect 1130 -47 1134 -43
rect 1278 -11 1282 -7
rect 1243 -36 1247 -32
rect 1379 -15 1383 -11
rect 1326 -36 1330 -32
rect 1296 -47 1300 -43
rect 1427 -30 1431 -26
rect 1397 -37 1401 -33
rect 1494 -15 1498 -11
rect 1476 -38 1480 -34
rect 1677 -19 1681 -15
rect 1542 -36 1546 -32
rect 1599 -35 1603 -31
rect 1635 -35 1639 -31
rect 1760 -18 1764 -14
rect 1725 -36 1729 -32
rect 1695 -47 1699 -43
rect 1861 -19 1865 -15
rect 1808 -36 1812 -32
rect 1843 -36 1847 -32
rect 1778 -47 1782 -43
rect 1891 -36 1895 -32
<< metal1 >>
rect -43 20 -39 24
rect -35 20 -28 24
rect -24 20 -17 24
rect -13 20 -3 24
rect 1 20 8 24
rect 12 20 19 24
rect 23 20 39 24
rect 43 20 53 24
rect 57 20 71 24
rect 75 20 87 24
rect 91 20 98 24
rect 102 20 109 24
rect 113 20 122 24
rect 126 20 136 24
rect 140 20 154 24
rect 158 20 170 24
rect 174 20 181 24
rect 185 20 192 24
rect 196 20 205 24
rect 209 20 219 24
rect 223 20 237 24
rect 241 20 253 24
rect 257 20 264 24
rect 268 20 275 24
rect 279 20 288 24
rect 292 20 302 24
rect 306 20 320 24
rect 324 20 336 24
rect 340 20 347 24
rect 351 20 358 24
rect 362 20 389 24
rect 393 20 403 24
rect 407 20 421 24
rect 425 20 437 24
rect 441 20 448 24
rect 452 20 459 24
rect 463 20 486 24
rect 490 20 500 24
rect 504 20 518 24
rect 522 20 552 24
rect 556 20 563 24
rect 567 20 574 24
rect 578 20 609 24
rect 613 20 620 24
rect 624 20 631 24
rect 635 20 645 24
rect 649 20 656 24
rect 660 20 667 24
rect 671 20 687 24
rect 691 20 701 24
rect 705 20 719 24
rect 723 20 735 24
rect 739 20 746 24
rect 750 20 757 24
rect 761 20 770 24
rect 774 20 784 24
rect 788 20 802 24
rect 806 20 818 24
rect 822 20 829 24
rect 833 20 840 24
rect 844 20 853 24
rect 857 20 867 24
rect 871 20 885 24
rect 889 20 901 24
rect 905 20 912 24
rect 916 20 923 24
rect 927 20 944 24
rect 948 20 955 24
rect 959 20 966 24
rect 970 20 980 24
rect 984 20 991 24
rect 995 20 1002 24
rect 1006 20 1022 24
rect 1026 20 1036 24
rect 1040 20 1054 24
rect 1058 20 1070 24
rect 1074 20 1081 24
rect 1085 20 1092 24
rect 1096 20 1105 24
rect 1109 20 1119 24
rect 1123 20 1137 24
rect 1141 20 1153 24
rect 1157 20 1164 24
rect 1168 20 1175 24
rect 1179 20 1188 24
rect 1192 20 1202 24
rect 1206 20 1220 24
rect 1224 20 1236 24
rect 1240 20 1247 24
rect 1251 20 1258 24
rect 1262 20 1271 24
rect 1275 20 1285 24
rect 1289 20 1303 24
rect 1307 20 1319 24
rect 1323 20 1330 24
rect 1334 20 1341 24
rect 1345 20 1372 24
rect 1376 20 1386 24
rect 1390 20 1404 24
rect 1408 20 1420 24
rect 1424 20 1431 24
rect 1435 20 1442 24
rect 1446 20 1469 24
rect 1473 20 1483 24
rect 1487 20 1501 24
rect 1505 20 1535 24
rect 1539 20 1546 24
rect 1550 20 1557 24
rect 1561 20 1592 24
rect 1596 20 1603 24
rect 1607 20 1614 24
rect 1618 20 1628 24
rect 1632 20 1639 24
rect 1643 20 1650 24
rect 1654 20 1670 24
rect 1674 20 1684 24
rect 1688 20 1702 24
rect 1706 20 1718 24
rect 1722 20 1729 24
rect 1733 20 1740 24
rect 1744 20 1753 24
rect 1757 20 1767 24
rect 1771 20 1785 24
rect 1789 20 1801 24
rect 1805 20 1812 24
rect 1816 20 1823 24
rect 1827 20 1836 24
rect 1840 20 1850 24
rect 1854 20 1868 24
rect 1872 20 1884 24
rect 1888 20 1895 24
rect 1899 20 1906 24
rect 1910 20 1913 24
rect -39 8 -35 20
rect -3 8 1 20
rect 39 8 43 20
rect 71 8 75 20
rect 87 8 91 20
rect 122 8 126 20
rect 154 8 158 20
rect 170 8 174 20
rect 205 8 209 20
rect 253 8 257 20
rect 288 8 292 20
rect 320 8 324 20
rect 336 8 340 20
rect 389 8 393 20
rect 421 8 425 20
rect 437 8 441 20
rect 486 8 490 20
rect 552 8 556 20
rect 609 8 613 20
rect 645 8 649 20
rect 687 8 691 20
rect 719 8 723 20
rect 735 8 739 20
rect 770 8 774 20
rect 802 8 806 20
rect 818 8 822 20
rect 853 8 857 20
rect 901 8 905 20
rect 944 8 948 20
rect 980 8 984 20
rect 1022 8 1026 20
rect 1054 8 1058 20
rect 1070 8 1074 20
rect 1105 8 1109 20
rect 1137 8 1141 20
rect 1153 8 1157 20
rect 1188 8 1192 20
rect 1236 8 1240 20
rect 1271 8 1275 20
rect 1303 8 1307 20
rect 1319 8 1323 20
rect 1372 8 1376 20
rect 1404 8 1408 20
rect 1420 8 1424 20
rect 1469 8 1473 20
rect 1535 8 1539 20
rect 1592 8 1596 20
rect 1628 8 1632 20
rect 1670 8 1674 20
rect 1702 8 1706 20
rect 1718 8 1722 20
rect 1753 8 1757 20
rect 1785 8 1789 20
rect 1801 8 1805 20
rect 1836 8 1840 20
rect 1884 8 1888 20
rect -38 -31 -34 -20
rect -21 -31 -17 0
rect -14 -31 -10 -29
rect 15 -31 19 0
rect 37 -19 46 -15
rect -38 -35 -32 -31
rect -21 -35 -10 -31
rect -6 -35 4 -31
rect 15 -35 38 -31
rect 53 -32 57 0
rect 105 -32 109 0
rect 114 -18 129 -14
rect 114 -23 118 -18
rect 136 -32 140 0
rect 188 -32 192 0
rect 204 -19 230 -15
rect 237 -32 241 0
rect 271 -32 275 0
rect 289 -11 295 -7
rect 282 -32 286 -22
rect 53 -35 94 -32
rect -48 -47 -39 -43
rect -21 -60 -17 -35
rect -6 -42 -2 -35
rect 15 -60 19 -35
rect 34 -43 38 -35
rect 71 -36 94 -35
rect 105 -36 115 -32
rect 34 -47 64 -43
rect 71 -60 75 -36
rect 105 -60 109 -36
rect 136 -35 177 -32
rect 154 -36 177 -35
rect 188 -36 212 -32
rect 219 -36 260 -32
rect 271 -36 286 -32
rect 302 -32 306 0
rect 354 -32 358 0
rect 376 -15 396 -11
rect 403 -26 407 0
rect 403 -30 444 -26
rect 302 -36 343 -32
rect 354 -36 375 -32
rect 116 -47 147 -43
rect 116 -50 120 -47
rect 154 -60 158 -36
rect 188 -60 192 -36
rect 219 -60 223 -36
rect 271 -60 275 -36
rect 282 -47 313 -43
rect 282 -50 286 -47
rect 320 -60 324 -36
rect 354 -60 358 -36
rect 371 -52 375 -36
rect 403 -37 405 -33
rect 410 -37 414 -33
rect 421 -60 425 -30
rect 455 -32 459 0
rect 464 -15 511 -11
rect 464 -32 468 -15
rect 518 -32 522 0
rect 570 -32 574 0
rect 610 -31 614 -24
rect 627 -31 631 0
rect 634 -31 638 -29
rect 663 -31 667 0
rect 685 -19 694 -15
rect 455 -36 468 -32
rect 455 -60 459 -36
rect 473 -38 493 -34
rect 500 -36 559 -32
rect 570 -36 588 -32
rect 610 -35 616 -31
rect 627 -35 638 -31
rect 642 -35 652 -31
rect 663 -35 686 -31
rect 701 -32 705 0
rect 753 -32 757 0
rect 762 -18 777 -14
rect 762 -23 766 -18
rect 784 -32 788 0
rect 836 -32 840 0
rect 852 -19 878 -15
rect 885 -32 889 0
rect 919 -32 923 0
rect 945 -31 949 -20
rect 962 -31 966 0
rect 969 -31 973 -29
rect 998 -31 1002 0
rect 1020 -19 1029 -15
rect 701 -35 742 -32
rect 473 -52 477 -38
rect 500 -60 504 -36
rect 570 -60 574 -36
rect 584 -52 588 -36
rect 605 -46 609 -42
rect 627 -60 631 -35
rect 642 -41 646 -35
rect 663 -60 667 -35
rect 682 -43 686 -35
rect 719 -36 742 -35
rect 753 -36 763 -32
rect 682 -47 712 -43
rect 719 -60 723 -36
rect 753 -60 757 -36
rect 784 -35 825 -32
rect 802 -36 825 -35
rect 836 -36 860 -32
rect 867 -36 908 -32
rect 919 -36 930 -32
rect 945 -35 951 -31
rect 962 -35 973 -31
rect 977 -35 987 -31
rect 998 -35 1021 -31
rect 1036 -32 1040 0
rect 1088 -32 1092 0
rect 1097 -18 1112 -14
rect 1097 -23 1101 -18
rect 1119 -32 1123 0
rect 1171 -32 1175 0
rect 1187 -19 1213 -15
rect 1220 -32 1224 0
rect 1254 -32 1258 0
rect 1272 -11 1278 -7
rect 1265 -32 1269 -22
rect 1036 -35 1077 -32
rect 764 -47 795 -43
rect 764 -50 768 -47
rect 802 -60 806 -36
rect 836 -60 840 -36
rect 867 -60 871 -36
rect 919 -60 923 -36
rect 935 -47 944 -43
rect 962 -60 966 -35
rect 977 -42 981 -35
rect 998 -60 1002 -35
rect 1017 -43 1021 -35
rect 1054 -36 1077 -35
rect 1088 -36 1098 -32
rect 1017 -47 1047 -43
rect 1054 -60 1058 -36
rect 1088 -60 1092 -36
rect 1119 -35 1160 -32
rect 1137 -36 1160 -35
rect 1171 -36 1195 -32
rect 1202 -36 1243 -32
rect 1254 -36 1269 -32
rect 1285 -32 1289 0
rect 1337 -32 1341 0
rect 1359 -15 1379 -11
rect 1386 -26 1390 0
rect 1386 -30 1427 -26
rect 1285 -36 1326 -32
rect 1337 -36 1358 -32
rect 1099 -47 1130 -43
rect 1099 -50 1103 -47
rect 1137 -60 1141 -36
rect 1171 -60 1175 -36
rect 1202 -60 1206 -36
rect 1254 -60 1258 -36
rect 1265 -47 1296 -43
rect 1265 -50 1269 -47
rect 1303 -60 1307 -36
rect 1337 -60 1341 -36
rect 1354 -52 1358 -36
rect 1363 -37 1388 -33
rect -39 -72 -35 -64
rect -3 -72 1 -64
rect 39 -72 43 -64
rect 87 -72 91 -64
rect 122 -72 126 -64
rect 170 -72 174 -64
rect 205 -72 209 -64
rect 237 -72 241 -64
rect 253 -72 257 -64
rect 288 -72 292 -64
rect 336 -72 340 -64
rect 389 -72 393 -64
rect 437 -72 441 -64
rect 486 -72 490 -64
rect 518 -72 522 -64
rect 552 -72 556 -64
rect 609 -72 613 -64
rect 645 -72 649 -64
rect 687 -72 691 -64
rect 735 -72 739 -64
rect 770 -72 774 -64
rect 818 -72 822 -64
rect 853 -72 857 -64
rect 885 -72 889 -64
rect 901 -72 905 -64
rect 944 -72 948 -64
rect 980 -72 984 -64
rect 1022 -72 1026 -64
rect 1070 -72 1074 -64
rect 1105 -72 1109 -64
rect 1153 -72 1157 -64
rect 1188 -72 1192 -64
rect 1220 -72 1224 -64
rect 1363 -63 1367 -37
rect 1393 -37 1397 -33
rect 1404 -60 1408 -30
rect 1438 -32 1442 0
rect 1447 -15 1494 -11
rect 1447 -32 1451 -15
rect 1501 -32 1505 0
rect 1553 -32 1557 0
rect 1593 -31 1597 -24
rect 1610 -31 1614 0
rect 1617 -31 1621 -29
rect 1646 -31 1650 0
rect 1668 -19 1677 -15
rect 1438 -36 1451 -32
rect 1438 -60 1442 -36
rect 1456 -38 1476 -34
rect 1483 -36 1542 -32
rect 1553 -36 1564 -32
rect 1593 -35 1599 -31
rect 1610 -35 1621 -31
rect 1625 -35 1635 -31
rect 1646 -35 1669 -31
rect 1684 -32 1688 0
rect 1736 -32 1740 0
rect 1745 -18 1760 -14
rect 1745 -23 1749 -18
rect 1767 -32 1771 0
rect 1819 -32 1823 0
rect 1835 -19 1861 -15
rect 1868 -32 1872 0
rect 1902 -32 1906 0
rect 1684 -35 1725 -32
rect 1456 -52 1460 -38
rect 1483 -60 1487 -36
rect 1553 -60 1557 -36
rect 1588 -46 1592 -42
rect 1610 -60 1614 -35
rect 1625 -41 1629 -35
rect 1646 -60 1650 -35
rect 1665 -43 1669 -35
rect 1702 -36 1725 -35
rect 1736 -36 1746 -32
rect 1665 -47 1695 -43
rect 1702 -60 1706 -36
rect 1736 -60 1740 -36
rect 1767 -35 1808 -32
rect 1785 -36 1808 -35
rect 1819 -36 1843 -32
rect 1850 -36 1891 -32
rect 1902 -36 1913 -32
rect 1747 -47 1778 -43
rect 1747 -50 1751 -47
rect 1785 -60 1789 -36
rect 1819 -60 1823 -36
rect 1850 -60 1854 -36
rect 1902 -60 1906 -36
rect 1236 -72 1240 -64
rect 1271 -72 1275 -64
rect 1319 -72 1323 -64
rect 1372 -72 1376 -64
rect 1420 -72 1424 -64
rect 1469 -72 1473 -64
rect 1501 -72 1505 -64
rect 1535 -72 1539 -64
rect 1592 -72 1596 -64
rect 1628 -72 1632 -64
rect 1670 -72 1674 -64
rect 1718 -72 1722 -64
rect 1753 -72 1757 -64
rect 1801 -72 1805 -64
rect 1836 -72 1840 -64
rect 1868 -72 1872 -64
rect 1884 -72 1888 -64
rect -43 -76 -39 -72
rect -35 -76 -25 -72
rect -21 -76 -14 -72
rect -10 -76 -3 -72
rect 1 -76 11 -72
rect 15 -76 22 -72
rect 26 -76 39 -72
rect 43 -76 53 -72
rect 57 -76 67 -72
rect 71 -76 87 -72
rect 91 -76 101 -72
rect 105 -76 112 -72
rect 116 -76 122 -72
rect 126 -76 136 -72
rect 140 -76 150 -72
rect 154 -76 170 -72
rect 174 -76 184 -72
rect 188 -76 195 -72
rect 199 -76 205 -72
rect 209 -76 219 -72
rect 223 -76 237 -72
rect 241 -76 253 -72
rect 257 -76 267 -72
rect 271 -76 278 -72
rect 282 -76 288 -72
rect 292 -76 302 -72
rect 306 -76 316 -72
rect 320 -76 336 -72
rect 340 -76 350 -72
rect 354 -76 361 -72
rect 365 -76 389 -72
rect 393 -76 403 -72
rect 407 -76 417 -72
rect 421 -76 437 -72
rect 441 -76 451 -72
rect 455 -76 462 -72
rect 466 -76 486 -72
rect 490 -76 500 -72
rect 504 -76 518 -72
rect 522 -76 552 -72
rect 556 -76 566 -72
rect 570 -76 577 -72
rect 581 -76 609 -72
rect 613 -76 623 -72
rect 627 -76 634 -72
rect 638 -76 645 -72
rect 649 -76 659 -72
rect 663 -76 670 -72
rect 674 -76 687 -72
rect 691 -76 701 -72
rect 705 -76 715 -72
rect 719 -76 735 -72
rect 739 -76 749 -72
rect 753 -76 760 -72
rect 764 -76 770 -72
rect 774 -76 784 -72
rect 788 -76 798 -72
rect 802 -76 818 -72
rect 822 -76 832 -72
rect 836 -76 843 -72
rect 847 -76 853 -72
rect 857 -76 867 -72
rect 871 -76 885 -72
rect 889 -76 901 -72
rect 905 -76 915 -72
rect 919 -76 926 -72
rect 930 -76 944 -72
rect 948 -76 958 -72
rect 962 -76 969 -72
rect 973 -76 980 -72
rect 984 -76 994 -72
rect 998 -76 1005 -72
rect 1009 -76 1022 -72
rect 1026 -76 1036 -72
rect 1040 -76 1050 -72
rect 1054 -76 1070 -72
rect 1074 -76 1084 -72
rect 1088 -76 1095 -72
rect 1099 -76 1105 -72
rect 1109 -76 1119 -72
rect 1123 -76 1133 -72
rect 1137 -76 1153 -72
rect 1157 -76 1167 -72
rect 1171 -76 1178 -72
rect 1182 -76 1188 -72
rect 1192 -76 1202 -72
rect 1206 -76 1220 -72
rect 1224 -76 1236 -72
rect 1240 -76 1250 -72
rect 1254 -76 1261 -72
rect 1265 -76 1271 -72
rect 1275 -76 1285 -72
rect 1289 -76 1299 -72
rect 1303 -76 1319 -72
rect 1323 -76 1333 -72
rect 1337 -76 1344 -72
rect 1348 -76 1372 -72
rect 1376 -76 1386 -72
rect 1390 -76 1400 -72
rect 1404 -76 1420 -72
rect 1424 -76 1434 -72
rect 1438 -76 1445 -72
rect 1449 -76 1469 -72
rect 1473 -76 1483 -72
rect 1487 -76 1501 -72
rect 1505 -76 1535 -72
rect 1539 -76 1549 -72
rect 1553 -76 1560 -72
rect 1564 -76 1592 -72
rect 1596 -76 1606 -72
rect 1610 -76 1617 -72
rect 1621 -76 1628 -72
rect 1632 -76 1642 -72
rect 1646 -76 1653 -72
rect 1657 -76 1670 -72
rect 1674 -76 1684 -72
rect 1688 -76 1698 -72
rect 1702 -76 1718 -72
rect 1722 -76 1732 -72
rect 1736 -76 1743 -72
rect 1747 -76 1753 -72
rect 1757 -76 1767 -72
rect 1771 -76 1781 -72
rect 1785 -76 1801 -72
rect 1805 -76 1815 -72
rect 1819 -76 1826 -72
rect 1830 -76 1836 -72
rect 1840 -76 1850 -72
rect 1854 -76 1868 -72
rect 1872 -76 1884 -72
rect 1888 -76 1898 -72
rect 1902 -76 1909 -72
<< m2contact >>
rect -38 -20 -33 -15
rect -14 -29 -9 -24
rect 32 -20 37 -15
rect 114 -28 119 -23
rect 199 -20 204 -15
rect 284 -12 289 -7
rect 282 -22 287 -17
rect -39 -47 -34 -42
rect -7 -47 -2 -42
rect 115 -37 120 -32
rect 371 -16 376 -11
rect 116 -55 121 -50
rect 282 -55 287 -50
rect 405 -38 410 -33
rect 371 -57 376 -52
rect 610 -24 615 -19
rect 634 -29 639 -24
rect 680 -20 685 -15
rect 762 -28 767 -23
rect 847 -20 852 -15
rect 945 -20 950 -15
rect 969 -29 974 -24
rect 1015 -20 1020 -15
rect 473 -57 478 -52
rect 600 -46 605 -41
rect 609 -46 614 -41
rect 584 -57 589 -52
rect 641 -46 646 -41
rect 763 -37 768 -32
rect 1097 -28 1102 -23
rect 1182 -20 1187 -15
rect 1267 -12 1272 -7
rect 1265 -22 1270 -17
rect 764 -55 769 -50
rect 944 -47 949 -42
rect 976 -47 981 -42
rect 1098 -37 1103 -32
rect 1354 -16 1359 -11
rect 1099 -55 1104 -50
rect 1265 -55 1270 -50
rect 1354 -57 1359 -52
rect 1388 -38 1393 -33
rect 1593 -24 1598 -19
rect 1617 -29 1622 -24
rect 1663 -20 1668 -15
rect 1745 -28 1750 -23
rect 1830 -20 1835 -15
rect 1456 -57 1461 -52
rect 1583 -46 1588 -41
rect 1592 -46 1597 -41
rect 1624 -46 1629 -41
rect 1746 -37 1751 -32
rect 1747 -55 1752 -50
rect 1362 -68 1367 -63
<< metal2 >>
rect -38 -11 284 -7
rect -38 -15 -34 -11
rect 945 -11 1267 -7
rect -33 -19 32 -15
rect 163 -19 199 -15
rect -9 -28 114 -24
rect 163 -32 167 -19
rect 945 -15 949 -11
rect 371 -17 375 -16
rect 287 -20 375 -17
rect 610 -19 680 -15
rect 287 -21 610 -20
rect 371 -24 610 -21
rect 811 -19 847 -15
rect 639 -28 762 -24
rect 811 -32 815 -19
rect 950 -19 1015 -15
rect 1146 -19 1182 -15
rect 974 -28 1097 -24
rect 1146 -32 1150 -19
rect 1354 -17 1358 -16
rect 1270 -20 1358 -17
rect 1593 -19 1663 -15
rect 1270 -21 1593 -20
rect 1354 -24 1593 -21
rect 1794 -19 1830 -15
rect 1622 -28 1745 -24
rect 1794 -32 1798 -19
rect 120 -36 167 -32
rect 768 -36 815 -32
rect 1103 -36 1150 -32
rect 1751 -36 1798 -32
rect 405 -42 409 -38
rect -34 -47 -7 -43
rect 405 -46 600 -42
rect 614 -46 641 -42
rect 1388 -42 1392 -38
rect -38 -51 -34 -47
rect -38 -55 116 -51
rect 121 -55 282 -51
rect 610 -51 614 -46
rect 949 -47 976 -43
rect 1388 -46 1583 -42
rect 1597 -46 1624 -42
rect 376 -57 473 -53
rect 610 -55 764 -51
rect 945 -51 949 -47
rect 945 -55 1099 -51
rect 1104 -55 1265 -51
rect 1593 -51 1597 -46
rect 1359 -57 1456 -53
rect 1593 -55 1747 -51
rect 1752 -55 1913 -51
rect 584 -85 588 -57
rect 1363 -85 1367 -68
rect 584 -89 1367 -85
<< labels >>
rlabel metal1 1561 -34 1561 -34 1 C2
rlabel metal1 1910 -35 1910 -35 7 S1
rlabel metal1 1367 -35 1367 -35 1 C1
rlabel metal1 946 -33 946 -33 1 A1
rlabel metal1 937 -45 937 -45 3 B1
rlabel metal1 1893 -74 1894 -73 1 GND
rlabel metal1 1846 -75 1847 -74 1 GND
rlabel metal1 1810 -74 1811 -73 1 GND
rlabel metal1 1764 -74 1765 -73 1 GND
rlabel metal1 1727 -74 1728 -73 1 GND
rlabel metal1 1680 -74 1681 -73 1 GND
rlabel metal1 1637 -75 1638 -74 1 GND
rlabel metal1 1600 -74 1601 -73 1 GND
rlabel metal1 1542 -74 1543 -73 1 GND
rlabel metal1 1477 -74 1478 -73 1 GND
rlabel metal1 1428 -75 1429 -74 1 GND
rlabel metal1 1327 -74 1328 -73 1 GND
rlabel metal1 1282 -74 1283 -73 1 GND
rlabel metal1 1245 -74 1246 -73 1 GND
rlabel metal1 1198 -74 1199 -73 1 GND
rlabel metal1 1427 22 1428 23 5 VDD
rlabel metal1 1478 22 1479 23 5 VDD
rlabel metal1 1542 22 1543 23 5 VDD
rlabel metal1 1600 21 1601 22 5 VDD
rlabel metal1 1637 22 1638 23 5 VDD
rlabel metal1 1677 22 1678 23 5 VDD
rlabel metal1 1725 22 1726 23 5 VDD
rlabel metal1 1762 21 1763 22 5 VDD
rlabel metal1 1809 22 1810 23 5 VDD
rlabel metal1 1845 21 1846 22 5 VDD
rlabel metal1 1892 22 1893 23 5 VDD
rlabel metal1 1327 22 1328 23 5 VDD
rlabel metal1 1282 22 1283 23 5 VDD
rlabel metal1 1244 22 1245 23 5 VDD
rlabel metal1 1198 22 1199 23 5 VDD
rlabel metal1 1383 -74 1383 -74 1 GND
rlabel metal1 1381 22 1381 22 5 VDD
rlabel metal1 1161 -75 1161 -75 1 GND
rlabel metal1 1115 -75 1115 -75 1 GND
rlabel metal1 1080 -73 1080 -73 1 GND
rlabel metal1 1033 -74 1033 -74 1 GND
rlabel metal1 989 -74 989 -74 1 GND
rlabel metal1 1162 22 1162 22 5 VDD
rlabel metal1 1077 22 1077 22 5 VDD
rlabel metal1 1115 22 1115 22 5 VDD
rlabel metal1 1033 22 1033 22 5 VDD
rlabel metal1 987 21 987 21 5 VDD
rlabel metal1 953 -74 953 -74 1 GND
rlabel metal1 951 22 951 22 5 VDD
rlabel metal1 404 -35 404 -35 1 Cin
rlabel metal1 910 -74 911 -73 1 GND
rlabel metal1 863 -75 864 -74 1 GND
rlabel metal1 827 -74 828 -73 1 GND
rlabel metal1 781 -74 782 -73 1 GND
rlabel metal1 744 -74 745 -73 1 GND
rlabel metal1 697 -74 698 -73 1 GND
rlabel metal1 654 -75 655 -74 1 GND
rlabel metal1 617 -74 618 -73 1 GND
rlabel metal1 559 -74 560 -73 1 GND
rlabel metal1 494 -74 495 -73 1 GND
rlabel metal1 445 -75 446 -74 1 GND
rlabel metal1 344 -74 345 -73 1 GND
rlabel metal1 299 -74 300 -73 1 GND
rlabel metal1 262 -74 263 -73 1 GND
rlabel metal1 215 -74 216 -73 1 GND
rlabel metal1 444 22 445 23 5 VDD
rlabel metal1 495 22 496 23 5 VDD
rlabel metal1 559 22 560 23 5 VDD
rlabel metal1 617 21 618 22 5 VDD
rlabel metal1 654 22 655 23 5 VDD
rlabel metal1 694 22 695 23 5 VDD
rlabel metal1 742 22 743 23 5 VDD
rlabel metal1 779 21 780 22 5 VDD
rlabel metal1 826 22 827 23 5 VDD
rlabel metal1 862 21 863 22 5 VDD
rlabel metal1 909 22 910 23 5 VDD
rlabel metal1 344 22 345 23 5 VDD
rlabel metal1 299 22 300 23 5 VDD
rlabel metal1 261 22 262 23 5 VDD
rlabel metal1 215 22 216 23 5 VDD
rlabel metal1 400 -74 400 -74 1 GND
rlabel metal1 398 22 398 22 5 VDD
rlabel metal1 178 -75 178 -75 1 GND
rlabel metal1 132 -75 132 -75 1 GND
rlabel metal1 97 -73 97 -73 1 GND
rlabel metal1 50 -74 50 -74 1 GND
rlabel metal1 6 -74 6 -74 1 GND
rlabel metal1 179 22 179 22 5 VDD
rlabel metal1 94 22 94 22 5 VDD
rlabel metal1 132 22 132 22 5 VDD
rlabel metal1 50 22 50 22 5 VDD
rlabel metal1 4 21 4 21 5 VDD
rlabel metal1 -30 -74 -30 -74 1 GND
rlabel metal1 -32 22 -32 22 5 VDD
rlabel metal1 578 -34 578 -34 1 C1
rlabel metal1 927 -34 927 -34 7 S0
rlabel metal1 -37 -33 -37 -33 1 A0
rlabel metal1 -47 -45 -47 -45 3 B0
<< end >>
