magic
tech scmos
timestamp 1730317458
<< nwell >>
rect -6 -6 28 14
<< ntransistor >>
rect 10 -64 12 -60
<< ptransistor >>
rect 10 0 12 8
<< ndiffusion >>
rect 4 -64 10 -60
rect 12 -64 18 -60
<< pdiffusion >>
rect 4 0 10 8
rect 12 0 18 8
<< ndcontact >>
rect 0 -64 4 -60
rect 18 -64 22 -60
<< pdcontact >>
rect 0 0 4 8
rect 18 0 22 8
<< psubstratepcontact >>
rect 0 -76 4 -72
rect 11 -76 15 -72
rect 22 -76 26 -72
<< nsubstratencontact >>
rect 0 20 4 24
rect 11 20 15 24
rect 22 20 26 24
<< polysilicon >>
rect 10 8 12 12
rect 10 -31 12 0
rect 11 -35 12 -31
rect 10 -60 12 -35
rect 10 -67 12 -64
<< polycontact >>
rect 7 -35 11 -31
<< metal1 >>
rect -4 20 0 24
rect 4 20 11 24
rect 15 20 22 24
rect 0 8 4 20
rect 18 -31 22 0
rect 3 -35 7 -31
rect 18 -35 27 -31
rect 18 -60 22 -35
rect 0 -72 4 -64
rect -4 -76 0 -72
rect 4 -76 11 -72
rect 15 -76 22 -72
<< labels >>
rlabel metal1 27 -35 27 -31 7 out
rlabel metal1 3 -35 3 -31 1 in
rlabel metal1 7 22 7 22 5 VDD
rlabel metal1 7 -74 7 -74 1 gnd
<< end >>
